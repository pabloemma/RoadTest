--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   11:41:00 03/01/2017
-- Design Name:   
-- Module Name:   C:/ML605/RoadTest_V2.02/decodeTB.vhd
-- Project Name:  RoadTest_V2.02
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: decode
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY decodeTB IS
END decodeTB;
 
ARCHITECTURE behavior OF decodeTB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT decode
    PORT(
         rst : IN  std_logic;
         clk : IN  std_logic;
         ena : IN  std_logic;
         hit_vector : IN  std_logic_vector(19 downto 0);
         quadrant : OUT  std_logic_vector(3 downto 0);
         sta1 : OUT  std_logic_vector(79 downto 0);
         sta2 : OUT  std_logic_vector(49 downto 0);
         sta4 : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal rst : std_logic := '0';
   signal clk : std_logic := '0';
   signal ena : std_logic := '0';
   signal hit_vector : std_logic_vector(19 downto 0) := (others => '0');

 	--Outputs
   signal quadrant : std_logic_vector(3 downto 0);
   signal sta1 : std_logic_vector(79 downto 0);
   signal sta2 : std_logic_vector(49 downto 0);
   signal sta4 : std_logic_vector(31 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: decode PORT MAP (
          rst => rst,
          clk => clk,
          ena => ena,
          hit_vector => hit_vector,
          quadrant => quadrant,
          sta1 => sta1,
          sta2 => sta2,
          sta4 => sta4
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 50 ns;	
		rst<='1';
		wait for 20 ns;
		rst<='0';
		
		wait for 30 ns;
		hit_vector<=B"1100_0010_0000_0110_0110";
		ena<='1';
		wait for 10 ns;
		hit_vector<=B"0000_0010_0000_0000_0000";
		ena<='0';

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
